library verilog;
use verilog.vl_types.all;
entity lab6problem3_vlg_vec_tst is
end lab6problem3_vlg_vec_tst;
