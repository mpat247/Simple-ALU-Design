library verilog;
use verilog.vl_types.all;
entity lab6problem2_vlg_vec_tst is
end lab6problem2_vlg_vec_tst;
